`include "./riscv_pkg.sv"
`include "./rvh_pkg.sv"
`include "./rvh_l1d_pkg.sv"
`include "./uop_encoding_pkg.sv"