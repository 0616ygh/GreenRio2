`ifndef __RISCV_PKG_SV__
`define __RISCV_PKG_SV__
`ifdef USE_VERILATOR
`include "rvh_pkg.sv"
`endif //USE_VERILATOR

package riscv_pkg;



endpackage

`endif