module tb_top;

//memory load





endmodule