`ifndef __RVH_PKG_SV__
`define __RVH_PKG_SV__

package rvh_pkg;


endpackage : rvh_pkg

`endif